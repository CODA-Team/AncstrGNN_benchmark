


.topckt INV i vdd vss zn
m1 zn i vss vss nch_lvt l=40e-9 w=155e-9 m=1 nf=1 
m0 zn i vdd vdd pch_lvt l=40e-9 w=205e-9 m=1 nf=1 
.ends INV
