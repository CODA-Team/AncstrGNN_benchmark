.topckt COMPARATOR_PRE_AMP clk crossn crossp gnd intern interp outm outp vdd _net0 _net1
xm0 gnd intern gnd gnd nch_lvt w=1.05e-6 l=1e-6 
xm22 gnd interp gnd gnd nch_lvt w=1.05e-6 l=1e-6 
xm16 outm crossp gnd gnd nch_lvt w=1.44e-6 l=40e-9 
xm17 outp crossn gnd gnd nch_lvt w=1.44e-6 l=40e-9 
xm4 crossn crossp intern gnd nch_lvt w=1.92e-6 l=40e-9 
xm3 crossp crossn interp gnd nch_lvt w=1.92e-6 l=40e-9 
xm7 net050 clk gnd gnd nch_lvt w=8.64e-6 l=40e-9 
xm5 intern _net0 net050 gnd nch_lvt w=9.6e-6 l=40e-9 
xm6 interp _net1 net050 gnd nch_lvt w=9.6e-6 l=40e-9 
xm8 outm crossp vdd vdd pch_lvt w=2.88e-6 l=40e-9 
xm18 intern clk vdd vdd pch_lvt w=1.92e-6 l=40e-9 
xm15 outp crossn vdd vdd pch_lvt w=2.88e-6 l=40e-9 
xm19 interp clk vdd vdd pch_lvt w=1.92e-6 l=40e-9 
xm10 crossn clk vdd vdd pch_lvt w=1.92e-6 l=40e-9 
xm12 crossp clk vdd vdd pch_lvt w=1.92e-6 l=40e-9 
xm14 crossn crossp vdd vdd pch_lvt w=3.84e-6 l=40e-9 
xm13 crossp crossn vdd vdd pch_lvt w=3.84e-6 l=40e-9 
.ends COMPARATOR_PRE_AMP

