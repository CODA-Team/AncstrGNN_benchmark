.topckt NRZ_TRI_DAC_v3_dnw dinn dinnb dinp dinpb ein einb gnd ioutn ioutp vbn1 vbn2 vbp1 vbp2 vcm vdddac
xm16 vbp2 vbp2 vbp2 vdddac pch w=4e-6 l=500e-9 
xm2 vcm2 vbp2 v2 vdddac pch w=4e-6 l=500e-9 
xm7 vcm einb vcm2 vdddac pch w=800e-9 l=40e-9 
xm17 ioutp dinnb vcm2 vdddac pch w=800e-9 l=40e-9 
xm6 ioutn dinpb vcm2 vdddac pch w=800e-9 l=40e-9 
xm3 v2 vbp1 vdddac vdddac pch w=6e-6 l=1.5e-6 
xm12 v1 vbn1 gnd gnd nch w=2.1e-6 l=1.5e-6 
xm13 vcm1 vbn2 v1 gnd nch w=4e-6 l=500e-9 
xm21 vbn2 vbn2 vbn2 gnd nch w=4e-6 l=500e-9 
xm18 ioutp dinp vcm1 gnd nch w=400e-9 l=40e-9 
xm15 ioutn dinn vcm1 gnd nch w=400e-9 l=40e-9 
xm14 vcm ein vcm1 gnd nch w=400e-9 l=40e-9 
.ends NRZ_TRI_DAC_v3_dnw

